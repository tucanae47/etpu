module dump();
    initial begin
        $dumpfile ("top_systolic.vcd");
        $dumpvars (0, top_systolic);
        #1;
    end
endmodule